
`timescale 1ns / 1ps
`include "Md5CoreTestMacros.v"


module Md5CoreTest();

reg clk, reset, test_all;
reg [31:0] count = 0;
reg [511:0] chunk;

wire [31:0] a, b, c, d;
wire [127:0] digest;

Md5Core uut (
  .clk(clk),
  .wordChunk(chunk),
  .A0('h67452301),
  .B0('hefcdab89),
  .C0('h98badcfe),
  .D0('h10325476),
  .A64(a),
  .B64(b),
  .C64(c),
  .D64(d),
  .digestValue(digest)
);

initial
  begin
    clk = 0;
    forever #2 clk = !clk;
  end

initial
  begin
    reset = 0;
    #5 reset = 1;
    #4 reset = 0;
  end

 //Test cases

 //"The quick brown fox jumps over the lazy dog."
`TestCase(
  1,
  test1,
  'hc209d9e4,
  'h1cfbd090,
  'hadff68a0,
  'hd0cb22df,
  'b00000000000000000000000000000000000000000000000000000001011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000010111001100111011011110110010000100000011110010111101001100001011011000010000001100101011010000111010000100000011100100110010101110110011011110010000001110011011100000110110101110101011010100010000001111000011011110110011000100000011011100111011101101111011100100110001000100000011010110110001101101001011101010111000100100000011001010110100001010100)

  //"The quick brown fox jumps over the lazy dog"
  `TestCase(
    2,
    test2,
    'h9d7d109e,
    'h82b62b37,
    'h351dd86b,
    'hd619a442,
    'b00000000000000000000000000000000000000000000000000000001010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001100111011011110110010000100000011110010111101001100001011011000010000001100101011010000111010000100000011100100110010101110110011011110010000001110011011100000110110101110101011010100010000001111000011011110110011000100000011011100111011101101111011100100110001000100000011010110110001101101001011101010111000100100000011001010110100001010100)

//"A"
`TestCase(
  3,
  test3,
  'h7062c57f,
  'ha80fa7e7,
  'hb735591a,
  'h29beac2e,
  'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000001000001)



//"Hello World"
`TestCase(
  4,
  test4,
  'h6f01aa92,
  'hfee76ce9,
  'h32f0ec6f,
  'h32a4df6c,
  'b00000000000000000000000000000000000000000000000000000000010110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000110010001101100011100100110111101010111001000000110111101101100011011000110010101001000)

//"
`TestCase(
  5,
  test5,
  'hd98c1dd4,
  'h04b2008f,
  'h980980e9,
  'h7e42f8ec,
  'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000)

`define Result test1&test2&test3&test4&test5

always @(posedge clk)  count <= count + 1;
always @(posedge clk)
       if(count == 71) test_all <= `Result;
endmodule

